module TOP();
	Vortex Vortex();
endmodule

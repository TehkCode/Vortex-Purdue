// Copyright © 2019-2023
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`include "VX_define.vh"

interface VX_schedule_if #(parameter WARP_CNT = `NUM_WARPS, parameter THREAD_CNT = `NUM_THREADS, parameter WARP_CNT_WIDTH = `LOG2UP(WARP_CNT)) ();

    typedef struct packed {
        logic [`UUID_WIDTH-1:0]     uuid;
        logic [WARP_CNT_WIDTH-1:0]       wid;
        logic [THREAD_CNT-1:0]    tmask;        
        logic [`XLEN-1:0]           PC;
    } data_t;

    logic  valid;
    data_t data;
    logic  ready;

    modport master (
        output valid,
        output data,
        input  ready
    );

    modport slave (
        input  valid,
        input  data,
        output ready
    );

endinterface
